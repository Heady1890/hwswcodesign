-------------------------------------------------------------------------------
-- Title      : D5m Camera
-- Project    : SPEAR - Scalable Processor for Embedded Applications in
--              Realtime Environment
-------------------------------------------------------------------------------
-- File       : ext_CamD5m.vhd
-- Author     : BSc Folie Simon
-- Company    : TU Wien - Institut fr technische Informatik
-- Created    : 2011-29-05
-- Last update: 2011-29-05
-- Platform   : Altera 
-------------------------------------------------------------------------------
-- Description:
--
-------------------------------------------------------------------------------


--------------------------------------------------------------------------------
-- LIBRARY
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.spear_pkg.all;
use work.pkg_camd5m_read.all;

architecture behaviour of ext_camd5m_read is
begin

end behaviour;




